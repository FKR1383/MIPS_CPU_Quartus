library verilog;
use verilog.vl_types.all;
entity Extender_vlg_vec_tst is
end Extender_vlg_vec_tst;
