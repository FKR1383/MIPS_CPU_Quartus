library verilog;
use verilog.vl_types.all;
entity InstructionMemory_vlg_vec_tst is
end InstructionMemory_vlg_vec_tst;
