library verilog;
use verilog.vl_types.all;
entity SCADDER_TEST is
    port(
        S               : out    vl_logic_vector(7 downto 0);
        CIN             : in     vl_logic;
        A               : in     vl_logic_vector(7 downto 0);
        B               : in     vl_logic_vector(7 downto 0)
    );
end SCADDER_TEST;
