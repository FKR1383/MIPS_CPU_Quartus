library verilog;
use verilog.vl_types.all;
entity FIFO_Branch_Predictor_vlg_vec_tst is
end FIFO_Branch_Predictor_vlg_vec_tst;
