library verilog;
use verilog.vl_types.all;
entity PIPE_vlg_vec_tst is
end PIPE_vlg_vec_tst;
