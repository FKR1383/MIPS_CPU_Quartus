library verilog;
use verilog.vl_types.all;
entity Practical3_vlg_vec_tst is
end Practical3_vlg_vec_tst;
