library verilog;
use verilog.vl_types.all;
entity SUB_8bit_vlg_vec_tst is
end SUB_8bit_vlg_vec_tst;
