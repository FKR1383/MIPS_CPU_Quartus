library verilog;
use verilog.vl_types.all;
entity OR8bit_vlg_vec_tst is
end OR8bit_vlg_vec_tst;
