library verilog;
use verilog.vl_types.all;
entity InstructionMemory_vlg_sample_tst is
    port(
        Address         : in     vl_logic_vector(7 downto 0);
        CLOCK           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end InstructionMemory_vlg_sample_tst;
