library verilog;
use verilog.vl_types.all;
entity Extender_vlg_check_tst is
    port(
        IMM_EXTEND      : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Extender_vlg_check_tst;
