library verilog;
use verilog.vl_types.all;
entity SCADDER_TEST_vlg_vec_tst is
end SCADDER_TEST_vlg_vec_tst;
