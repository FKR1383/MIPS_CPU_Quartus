library verilog;
use verilog.vl_types.all;
entity Control_Multi_Cycle_vlg_vec_tst is
end Control_Multi_Cycle_vlg_vec_tst;
