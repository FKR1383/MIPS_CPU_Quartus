library verilog;
use verilog.vl_types.all;
entity PIPE1_Negedge_vlg_vec_tst is
end PIPE1_Negedge_vlg_vec_tst;
