library verilog;
use verilog.vl_types.all;
entity FLUSH_UNIT_vlg_vec_tst is
end FLUSH_UNIT_vlg_vec_tst;
