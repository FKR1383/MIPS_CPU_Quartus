library verilog;
use verilog.vl_types.all;
entity MIPS_CPU_vlg_vec_tst is
end MIPS_CPU_vlg_vec_tst;
