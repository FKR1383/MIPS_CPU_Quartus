library verilog;
use verilog.vl_types.all;
entity MIPS_CPU_MULTI_CYCLE_vlg_sample_tst is
    port(
        CLOCK           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end MIPS_CPU_MULTI_CYCLE_vlg_sample_tst;
