library verilog;
use verilog.vl_types.all;
entity Booth_Multiplier_vlg_vec_tst is
end Booth_Multiplier_vlg_vec_tst;
